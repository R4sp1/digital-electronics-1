------------------------------------------------------------
--
-- Example of 2-bit binary comparator using the when/else
-- assignments.
-- EDA Playground
--
-- Copyright (c) 2020-Present Tomas Fryza
-- Dept. of Radio Electronics, Brno Univ. of Technology, Czechia
-- This work is licensed under the terms of the MIT license.
--
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

------------------------------------------------------------
-- Entity declaration for 2-bit binary comparator
------------------------------------------------------------
entity comparator_2bit is
    port(
        b_i           : in  std_logic_vector(2 - 1 downto 0);	--DATA B
        a_i           : in	std_logic_vector(2 - 1 downto 0);	--DATA A
        B_greater_A_o : out	std_logic;							--B is greater then A
        B_equals_A_o  : out	std_logic;							--B equals A
        B_less_A_o    : out std_logic  							--B is less than A
    );
end entity comparator_2bit;

------------------------------------------------------------
-- Architecture body for 2-bit binary comparator
------------------------------------------------------------
architecture Behavioral of comparator_2bit is
begin
    B_greater_A_o <= '1' when (b_i > a_i) else '0';
    B_equals_A_o  <= '1' when (b_i = a_i) else '0';
    B_less_A_o    <= '1' when (b_i < a_i) else '0';

end architecture Behavioral;
